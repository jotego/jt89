/*  This file is part of JT89.

    JT89 is free software: you can redistribute it and/or modify
    it under the terms of the GNU General Public License as published by
    the Free Software Foundation, either version 3 of the License, or
    (at your option) any later version.

    JT89 is distributed in the hope that it will be useful,
    but WITHOUT ANY WARRANTY; without even the implied warranty of
    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
    GNU General Public License for more details.

    You should have received a copy of the GNU General Public License
    along with JT89.  If not, see <http://www.gnu.org/licenses/>.

    Author: Jose Tejada Gomez. Twitter: @topapate
    Version: 1.0
    Date: December, 1st 2018
   
    */

module jt89_mixer #(parameter bw=9)(
    input            rst,
    input            clk,
    input            clk_en,
    input            cen_16,
    input     [bw-1:0] ch0,
    input     [bw-1:0] ch1,
    input     [bw-1:0] ch2,
    input     [bw-1:0] noise,
    output    [bw+1:0] sound
);

reg signed [bw+1:0] fresh, old;

always @(*)
    fresh = 
        {2'b0, ch0   }+
        {2'b0, ch1   }+
        {2'b0, ch2   }+
        {2'b0, noise };

// Comb filter
localparam fbw=bw+7; // filter bit width
reg signed [fbw-1:0] comb1, old_comb1, comb2;
always @(posedge clk) if(cen_16) begin
    old <= fresh;
    comb1 <= {{(fbw-bw-2){1'b0}},fresh}-{{(fbw-bw-2){1'b0}},old};
    old_comb1 <= comb1;
    comb2 <= comb1-old_comb1;
end

// interpolator x16
reg signed [fbw-1:0] interp;
always @(posedge clk) if(clk_en) // clk_en = 16xcen_16
    interp <= cen_16 ? comb2 : {fbw{1'b0}};

// integrator
reg signed [fbw-1:0] integ1, integ2;
always @(posedge clk) 
    if( rst ) begin
        integ1 <= {fbw{1'b0}};
        integ2 <= {fbw{1'b0}};
    end else if(clk_en) begin
        integ1 <= integ1 + interp;
        integ2 <= integ2 + integ1;
    end
// scale back
assign sound = integ2[fbw-1] ? {bw+2{1'b0}} : // limit at zero
     integ2[fbw-2:fbw-bw-3]; // drop the sign bit

endmodule